/* String Descriptors */
localparam BOARD_VID = 16'h1d50;
localparam BOARD_PID = 16'h615d;
localparam BOARD_MFR_NAME = "oskirby";
localparam BOARD_PRODUCT_NAME = "Logicbone ECP5";
localparam BOARD_SERIAL = "123456";
